entity tb is
end entity;

architecture rg2 of tb is
begin
  process is

  begin

  end process;
end architecture;

